module EXE_Stage (
  input         clk,
  input         rst,
  input [31:0]  pc_in,
  output [31:0] pc
  );

endmodule
