module ConditionCheck (
  input [3:0]   cond,
  input [3:0]   sr,
  
  output        result
  );

endmodule

