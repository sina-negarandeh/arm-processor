module ID_Stage_Reg (
  input             clk,
  input             rst,
  output [31:0]     pc_in,
  output reg [31:0] pc
  );

endmodule
